// Nios2.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module Nios2 (
		output wire        audio_clk_clk,             //           audio_clk.clk
		input  wire        audio_pll_ref_clk_clk,     //   audio_pll_ref_clk.clk
		input  wire        audio_pll_ref_reset_reset, // audio_pll_ref_reset.reset
		input  wire        audiocore_ADCDAT,          //           audiocore.ADCDAT
		input  wire        audiocore_ADCLRCK,         //                    .ADCLRCK
		input  wire        audiocore_BCLK,            //                    .BCLK
		output wire        audiocore_DACDAT,          //                    .DACDAT
		input  wire        audiocore_DACLRCK,         //                    .DACLRCK
		inout  wire        avconfig_SDAT,             //            avconfig.SDAT
		output wire        avconfig_SCLK,             //                    .SCLK
		input  wire        clk_clk,                   //                 clk.clk
		inout  wire [31:0] gpio_expansion_export,     //      gpio_expansion.export
		output wire [6:0]  hex0_export,               //                hex0.export
		output wire [6:0]  hex1_export,               //                hex1.export
		output wire [6:0]  hex2_export,               //                hex2.export
		output wire [6:0]  hex3_export,               //                hex3.export
		output wire [6:0]  hex4_export,               //                hex4.export
		output wire [6:0]  hex5_export,               //                hex5.export
		output wire [6:0]  hex6_export,               //                hex6.export
		output wire [6:0]  hex7_export,               //                hex7.export
		input  wire [3:0]  keys_export,               //                keys.export
		output wire [7:0]  ledg_export,               //                ledg.export
		output wire [17:0] ledr_export,               //                ledr.export
		input  wire        reset_reset,               //               reset.reset
		output wire        sdram_clk_clk,             //           sdram_clk.clk
		output wire [12:0] sdram_wire_addr,           //          sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,             //                    .ba
		output wire        sdram_wire_cas_n,          //                    .cas_n
		output wire        sdram_wire_cke,            //                    .cke
		output wire        sdram_wire_cs_n,           //                    .cs_n
		inout  wire [31:0] sdram_wire_dq,             //                    .dq
		output wire [3:0]  sdram_wire_dqm,            //                    .dqm
		output wire        sdram_wire_ras_n,          //                    .ras_n
		output wire        sdram_wire_we_n,           //                    .we_n
		input  wire [17:0] switches_export            //            switches.export
	);

	wire         clocks_sys_clk_clk;                                                            // clocks:sys_clk_clk -> [AudioCore:clk, GPIO_Expansion:clk, HEX0:clk, HEX1:clk, HEX2:clk, HEX3:clk, HEX4:clk, HEX5:clk, HEX6:clk, HEX7:clk, KEYs:clk, LEDG:clk, LEDR:clk, audio_and_video_config_0:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:clocks_sys_clk_clk, myCPU:clk, rst_controller:clk, sdram:clk, switches:clk, sysid_qsys_0:clock, timer0:clk]
	wire  [31:0] mycpu_data_master_readdata;                                                    // mm_interconnect_0:myCPU_data_master_readdata -> myCPU:d_readdata
	wire         mycpu_data_master_waitrequest;                                                 // mm_interconnect_0:myCPU_data_master_waitrequest -> myCPU:d_waitrequest
	wire         mycpu_data_master_debugaccess;                                                 // myCPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:myCPU_data_master_debugaccess
	wire  [27:0] mycpu_data_master_address;                                                     // myCPU:d_address -> mm_interconnect_0:myCPU_data_master_address
	wire   [3:0] mycpu_data_master_byteenable;                                                  // myCPU:d_byteenable -> mm_interconnect_0:myCPU_data_master_byteenable
	wire         mycpu_data_master_read;                                                        // myCPU:d_read -> mm_interconnect_0:myCPU_data_master_read
	wire         mycpu_data_master_readdatavalid;                                               // mm_interconnect_0:myCPU_data_master_readdatavalid -> myCPU:d_readdatavalid
	wire         mycpu_data_master_write;                                                       // myCPU:d_write -> mm_interconnect_0:myCPU_data_master_write
	wire  [31:0] mycpu_data_master_writedata;                                                   // myCPU:d_writedata -> mm_interconnect_0:myCPU_data_master_writedata
	wire  [31:0] mycpu_instruction_master_readdata;                                             // mm_interconnect_0:myCPU_instruction_master_readdata -> myCPU:i_readdata
	wire         mycpu_instruction_master_waitrequest;                                          // mm_interconnect_0:myCPU_instruction_master_waitrequest -> myCPU:i_waitrequest
	wire  [27:0] mycpu_instruction_master_address;                                              // myCPU:i_address -> mm_interconnect_0:myCPU_instruction_master_address
	wire         mycpu_instruction_master_read;                                                 // myCPU:i_read -> mm_interconnect_0:myCPU_instruction_master_read
	wire         mycpu_instruction_master_readdatavalid;                                        // mm_interconnect_0:myCPU_instruction_master_readdatavalid -> myCPU:i_readdatavalid
	wire         mm_interconnect_0_audiocore_avalon_audio_slave_chipselect;                     // mm_interconnect_0:AudioCore_avalon_audio_slave_chipselect -> AudioCore:chipselect
	wire  [31:0] mm_interconnect_0_audiocore_avalon_audio_slave_readdata;                       // AudioCore:readdata -> mm_interconnect_0:AudioCore_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audiocore_avalon_audio_slave_address;                        // mm_interconnect_0:AudioCore_avalon_audio_slave_address -> AudioCore:address
	wire         mm_interconnect_0_audiocore_avalon_audio_slave_read;                           // mm_interconnect_0:AudioCore_avalon_audio_slave_read -> AudioCore:read
	wire         mm_interconnect_0_audiocore_avalon_audio_slave_write;                          // mm_interconnect_0:AudioCore_avalon_audio_slave_write -> AudioCore:write
	wire  [31:0] mm_interconnect_0_audiocore_avalon_audio_slave_writedata;                      // mm_interconnect_0:AudioCore_avalon_audio_slave_writedata -> AudioCore:writedata
	wire  [31:0] mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata;    // audio_and_video_config_0:readdata -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest; // audio_and_video_config_0:waitrequest -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address;     // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_address -> audio_and_video_config_0:address
	wire         mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read;        // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_read -> audio_and_video_config_0:read
	wire   [3:0] mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable;  // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_byteenable -> audio_and_video_config_0:byteenable
	wire         mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write;       // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_write -> audio_and_video_config_0:write
	wire  [31:0] mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata;   // mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_writedata -> audio_and_video_config_0:writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                      // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                   // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                         // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                          // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_mycpu_jtag_debug_module_readdata;                            // myCPU:jtag_debug_module_readdata -> mm_interconnect_0:myCPU_jtag_debug_module_readdata
	wire         mm_interconnect_0_mycpu_jtag_debug_module_waitrequest;                         // myCPU:jtag_debug_module_waitrequest -> mm_interconnect_0:myCPU_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_mycpu_jtag_debug_module_debugaccess;                         // mm_interconnect_0:myCPU_jtag_debug_module_debugaccess -> myCPU:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_mycpu_jtag_debug_module_address;                             // mm_interconnect_0:myCPU_jtag_debug_module_address -> myCPU:jtag_debug_module_address
	wire         mm_interconnect_0_mycpu_jtag_debug_module_read;                                // mm_interconnect_0:myCPU_jtag_debug_module_read -> myCPU:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_mycpu_jtag_debug_module_byteenable;                          // mm_interconnect_0:myCPU_jtag_debug_module_byteenable -> myCPU:jtag_debug_module_byteenable
	wire         mm_interconnect_0_mycpu_jtag_debug_module_write;                               // mm_interconnect_0:myCPU_jtag_debug_module_write -> myCPU:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_mycpu_jtag_debug_module_writedata;                           // mm_interconnect_0:myCPU_jtag_debug_module_writedata -> myCPU:jtag_debug_module_writedata
	wire         mm_interconnect_0_ledr_s1_chipselect;                                          // mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                                            // LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                                             // mm_interconnect_0:LEDR_s1_address -> LEDR:address
	wire         mm_interconnect_0_ledr_s1_write;                                               // mm_interconnect_0:LEDR_s1_write -> LEDR:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                                           // mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	wire         mm_interconnect_0_keys_s1_chipselect;                                          // mm_interconnect_0:KEYs_s1_chipselect -> KEYs:chipselect
	wire  [31:0] mm_interconnect_0_keys_s1_readdata;                                            // KEYs:readdata -> mm_interconnect_0:KEYs_s1_readdata
	wire   [1:0] mm_interconnect_0_keys_s1_address;                                             // mm_interconnect_0:KEYs_s1_address -> KEYs:address
	wire         mm_interconnect_0_keys_s1_write;                                               // mm_interconnect_0:KEYs_s1_write -> KEYs:write_n
	wire  [31:0] mm_interconnect_0_keys_s1_writedata;                                           // mm_interconnect_0:KEYs_s1_writedata -> KEYs:writedata
	wire         mm_interconnect_0_switches_s1_chipselect;                                      // mm_interconnect_0:switches_s1_chipselect -> switches:chipselect
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                                        // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                                         // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_switches_s1_write;                                           // mm_interconnect_0:switches_s1_write -> switches:write_n
	wire  [31:0] mm_interconnect_0_switches_s1_writedata;                                       // mm_interconnect_0:switches_s1_writedata -> switches:writedata
	wire         mm_interconnect_0_ledg_s1_chipselect;                                          // mm_interconnect_0:LEDG_s1_chipselect -> LEDG:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                                            // LEDG:readdata -> mm_interconnect_0:LEDG_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                                             // mm_interconnect_0:LEDG_s1_address -> LEDG:address
	wire         mm_interconnect_0_ledg_s1_write;                                               // mm_interconnect_0:LEDG_s1_write -> LEDG:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                                           // mm_interconnect_0:LEDG_s1_writedata -> LEDG:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                         // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                           // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                        // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                            // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                               // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                                         // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                      // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                              // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                                          // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_hex0_s1_chipselect;                                          // mm_interconnect_0:HEX0_s1_chipselect -> HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex0_s1_readdata;                                            // HEX0:readdata -> mm_interconnect_0:HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_s1_address;                                             // mm_interconnect_0:HEX0_s1_address -> HEX0:address
	wire         mm_interconnect_0_hex0_s1_write;                                               // mm_interconnect_0:HEX0_s1_write -> HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex0_s1_writedata;                                           // mm_interconnect_0:HEX0_s1_writedata -> HEX0:writedata
	wire         mm_interconnect_0_hex1_s1_chipselect;                                          // mm_interconnect_0:HEX1_s1_chipselect -> HEX1:chipselect
	wire  [31:0] mm_interconnect_0_hex1_s1_readdata;                                            // HEX1:readdata -> mm_interconnect_0:HEX1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex1_s1_address;                                             // mm_interconnect_0:HEX1_s1_address -> HEX1:address
	wire         mm_interconnect_0_hex1_s1_write;                                               // mm_interconnect_0:HEX1_s1_write -> HEX1:write_n
	wire  [31:0] mm_interconnect_0_hex1_s1_writedata;                                           // mm_interconnect_0:HEX1_s1_writedata -> HEX1:writedata
	wire         mm_interconnect_0_hex2_s1_chipselect;                                          // mm_interconnect_0:HEX2_s1_chipselect -> HEX2:chipselect
	wire  [31:0] mm_interconnect_0_hex2_s1_readdata;                                            // HEX2:readdata -> mm_interconnect_0:HEX2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex2_s1_address;                                             // mm_interconnect_0:HEX2_s1_address -> HEX2:address
	wire         mm_interconnect_0_hex2_s1_write;                                               // mm_interconnect_0:HEX2_s1_write -> HEX2:write_n
	wire  [31:0] mm_interconnect_0_hex2_s1_writedata;                                           // mm_interconnect_0:HEX2_s1_writedata -> HEX2:writedata
	wire         mm_interconnect_0_hex3_s1_chipselect;                                          // mm_interconnect_0:HEX3_s1_chipselect -> HEX3:chipselect
	wire  [31:0] mm_interconnect_0_hex3_s1_readdata;                                            // HEX3:readdata -> mm_interconnect_0:HEX3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_s1_address;                                             // mm_interconnect_0:HEX3_s1_address -> HEX3:address
	wire         mm_interconnect_0_hex3_s1_write;                                               // mm_interconnect_0:HEX3_s1_write -> HEX3:write_n
	wire  [31:0] mm_interconnect_0_hex3_s1_writedata;                                           // mm_interconnect_0:HEX3_s1_writedata -> HEX3:writedata
	wire         mm_interconnect_0_hex4_s1_chipselect;                                          // mm_interconnect_0:HEX4_s1_chipselect -> HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex4_s1_readdata;                                            // HEX4:readdata -> mm_interconnect_0:HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex4_s1_address;                                             // mm_interconnect_0:HEX4_s1_address -> HEX4:address
	wire         mm_interconnect_0_hex4_s1_write;                                               // mm_interconnect_0:HEX4_s1_write -> HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex4_s1_writedata;                                           // mm_interconnect_0:HEX4_s1_writedata -> HEX4:writedata
	wire         mm_interconnect_0_hex5_s1_chipselect;                                          // mm_interconnect_0:HEX5_s1_chipselect -> HEX5:chipselect
	wire  [31:0] mm_interconnect_0_hex5_s1_readdata;                                            // HEX5:readdata -> mm_interconnect_0:HEX5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_s1_address;                                             // mm_interconnect_0:HEX5_s1_address -> HEX5:address
	wire         mm_interconnect_0_hex5_s1_write;                                               // mm_interconnect_0:HEX5_s1_write -> HEX5:write_n
	wire  [31:0] mm_interconnect_0_hex5_s1_writedata;                                           // mm_interconnect_0:HEX5_s1_writedata -> HEX5:writedata
	wire         mm_interconnect_0_hex6_s1_chipselect;                                          // mm_interconnect_0:HEX6_s1_chipselect -> HEX6:chipselect
	wire  [31:0] mm_interconnect_0_hex6_s1_readdata;                                            // HEX6:readdata -> mm_interconnect_0:HEX6_s1_readdata
	wire   [1:0] mm_interconnect_0_hex6_s1_address;                                             // mm_interconnect_0:HEX6_s1_address -> HEX6:address
	wire         mm_interconnect_0_hex6_s1_write;                                               // mm_interconnect_0:HEX6_s1_write -> HEX6:write_n
	wire  [31:0] mm_interconnect_0_hex6_s1_writedata;                                           // mm_interconnect_0:HEX6_s1_writedata -> HEX6:writedata
	wire         mm_interconnect_0_hex7_s1_chipselect;                                          // mm_interconnect_0:HEX7_s1_chipselect -> HEX7:chipselect
	wire  [31:0] mm_interconnect_0_hex7_s1_readdata;                                            // HEX7:readdata -> mm_interconnect_0:HEX7_s1_readdata
	wire   [1:0] mm_interconnect_0_hex7_s1_address;                                             // mm_interconnect_0:HEX7_s1_address -> HEX7:address
	wire         mm_interconnect_0_hex7_s1_write;                                               // mm_interconnect_0:HEX7_s1_write -> HEX7:write_n
	wire  [31:0] mm_interconnect_0_hex7_s1_writedata;                                           // mm_interconnect_0:HEX7_s1_writedata -> HEX7:writedata
	wire         mm_interconnect_0_timer0_s1_chipselect;                                        // mm_interconnect_0:timer0_s1_chipselect -> timer0:chipselect
	wire  [15:0] mm_interconnect_0_timer0_s1_readdata;                                          // timer0:readdata -> mm_interconnect_0:timer0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer0_s1_address;                                           // mm_interconnect_0:timer0_s1_address -> timer0:address
	wire         mm_interconnect_0_timer0_s1_write;                                             // mm_interconnect_0:timer0_s1_write -> timer0:write_n
	wire  [15:0] mm_interconnect_0_timer0_s1_writedata;                                         // mm_interconnect_0:timer0_s1_writedata -> timer0:writedata
	wire         mm_interconnect_0_gpio_expansion_s1_chipselect;                                // mm_interconnect_0:GPIO_Expansion_s1_chipselect -> GPIO_Expansion:chipselect
	wire  [31:0] mm_interconnect_0_gpio_expansion_s1_readdata;                                  // GPIO_Expansion:readdata -> mm_interconnect_0:GPIO_Expansion_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_expansion_s1_address;                                   // mm_interconnect_0:GPIO_Expansion_s1_address -> GPIO_Expansion:address
	wire         mm_interconnect_0_gpio_expansion_s1_write;                                     // mm_interconnect_0:GPIO_Expansion_s1_write -> GPIO_Expansion:write_n
	wire  [31:0] mm_interconnect_0_gpio_expansion_s1_writedata;                                 // mm_interconnect_0:GPIO_Expansion_s1_writedata -> GPIO_Expansion:writedata
	wire         irq_mapper_receiver0_irq;                                                      // AudioCore:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                      // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                      // timer0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                      // KEYs:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                      // GPIO_Expansion:irq -> irq_mapper:receiver4_irq
	wire  [31:0] mycpu_d_irq_irq;                                                               // irq_mapper:sender_irq -> myCPU:d_irq
	wire         rst_controller_reset_out_reset;                                                // rst_controller:reset_out -> [AudioCore:reset, GPIO_Expansion:reset_n, HEX0:reset_n, HEX1:reset_n, HEX2:reset_n, HEX3:reset_n, HEX4:reset_n, HEX5:reset_n, HEX6:reset_n, HEX7:reset_n, KEYs:reset_n, LEDG:reset_n, LEDR:reset_n, audio_and_video_config_0:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:myCPU_reset_n_reset_bridge_in_reset_reset, myCPU:reset_n, rst_translator:in_reset, sdram:reset_n, switches:reset_n, sysid_qsys_0:reset_n, timer0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                            // rst_controller:reset_req -> [myCPU:reset_req, rst_translator:reset_req_in]
	wire         mycpu_jtag_debug_module_reset_reset;                                           // myCPU:jtag_debug_module_resetrequest -> rst_controller:reset_in0
	wire         clocks_reset_source_reset;                                                     // clocks:reset_source_reset -> rst_controller:reset_in1

	Nios2_AudioCore audiocore (
		.clk         (clocks_sys_clk_clk),                                        //                clk.clk
		.reset       (rst_controller_reset_out_reset),                            //              reset.reset
		.address     (mm_interconnect_0_audiocore_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audiocore_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audiocore_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audiocore_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audiocore_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audiocore_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver0_irq),                                  //          interrupt.irq
		.AUD_ADCDAT  (audiocore_ADCDAT),                                          // external_interface.export
		.AUD_ADCLRCK (audiocore_ADCLRCK),                                         //                   .export
		.AUD_BCLK    (audiocore_BCLK),                                            //                   .export
		.AUD_DACDAT  (audiocore_DACDAT),                                          //                   .export
		.AUD_DACLRCK (audiocore_DACLRCK)                                          //                   .export
	);

	Nios2_GPIO_Expansion gpio_expansion (
		.clk        (clocks_sys_clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_gpio_expansion_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_expansion_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_expansion_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_expansion_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_expansion_s1_readdata),   //                    .readdata
		.bidir_port (gpio_expansion_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                        //                 irq.irq
	);

	Nios2_HEX0 hex0 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex0_export)                           // external_connection.export
	);

	Nios2_HEX0 hex1 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex1_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                           // external_connection.export
	);

	Nios2_HEX0 hex2 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex2_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                           // external_connection.export
	);

	Nios2_HEX0 hex3 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_s1_readdata),   //                    .readdata
		.out_port   (hex3_export)                           // external_connection.export
	);

	Nios2_HEX0 hex4 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex4_export)                           // external_connection.export
	);

	Nios2_HEX0 hex5 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_s1_readdata),   //                    .readdata
		.out_port   (hex5_export)                           // external_connection.export
	);

	Nios2_HEX0 hex6 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex6_s1_readdata),   //                    .readdata
		.out_port   (hex6_export)                           // external_connection.export
	);

	Nios2_HEX0 hex7 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex7_s1_readdata),   //                    .readdata
		.out_port   (hex7_export)                           // external_connection.export
	);

	Nios2_KEYs keys (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_keys_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keys_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keys_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keys_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keys_s1_readdata),   //                    .readdata
		.in_port    (keys_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)              //                 irq.irq
	);

	Nios2_LEDG ledg (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                           // external_connection.export
	);

	Nios2_LEDR ledr (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	Nios2_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (clocks_sys_clk_clk),                                                            //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                                //                  reset.reset
		.address     (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (avconfig_SDAT),                                                                 //     external_interface.export
		.I2C_SCLK    (avconfig_SCLK)                                                                  //                       .export
	);

	Nios2_audio_pll_0 audio_pll_0 (
		.ref_clk_clk        (audio_pll_ref_clk_clk),     //      ref_clk.clk
		.ref_reset_reset    (audio_pll_ref_reset_reset), //    ref_reset.reset
		.audio_clk_clk      (audio_clk_clk),             //    audio_clk.clk
		.reset_source_reset ()                           // reset_source.reset
	);

	Nios2_clocks clocks (
		.ref_clk_clk        (clk_clk),                   //      ref_clk.clk
		.ref_reset_reset    (reset_reset),               //    ref_reset.reset
		.sys_clk_clk        (clocks_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),             //    sdram_clk.clk
		.reset_source_reset (clocks_reset_source_reset)  // reset_source.reset
	);

	Nios2_jtag_uart_0 jtag_uart_0 (
		.clk            (clocks_sys_clk_clk),                                          //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	Nios2_myCPU mycpu (
		.clk                                   (clocks_sys_clk_clk),                                    //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (mycpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (mycpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (mycpu_data_master_read),                                //                          .read
		.d_readdata                            (mycpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (mycpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (mycpu_data_master_write),                               //                          .write
		.d_writedata                           (mycpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (mycpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (mycpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (mycpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (mycpu_instruction_master_read),                         //                          .read
		.i_readdata                            (mycpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (mycpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (mycpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (mycpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (mycpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_mycpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_mycpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_mycpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_mycpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_mycpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_mycpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_mycpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_mycpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	Nios2_sdram sdram (
		.clk            (clocks_sys_clk_clk),                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	Nios2_switches switches (
		.clk        (clocks_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_switches_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_switches_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_switches_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_switches_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_switches_s1_readdata),   //                    .readdata
		.in_port    (switches_export)                           // external_connection.export
	);

	Nios2_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clocks_sys_clk_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	Nios2_timer0 timer0 (
		.clk        (clocks_sys_clk_clk),                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_0_timer0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                //   irq.irq
	);

	Nios2_mm_interconnect_0 mm_interconnect_0 (
		.clocks_sys_clk_clk                                          (clocks_sys_clk_clk),                                                            //                                  clocks_sys_clk.clk
		.myCPU_reset_n_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                                                //             myCPU_reset_n_reset_bridge_in_reset.reset
		.myCPU_data_master_address                                   (mycpu_data_master_address),                                                     //                               myCPU_data_master.address
		.myCPU_data_master_waitrequest                               (mycpu_data_master_waitrequest),                                                 //                                                .waitrequest
		.myCPU_data_master_byteenable                                (mycpu_data_master_byteenable),                                                  //                                                .byteenable
		.myCPU_data_master_read                                      (mycpu_data_master_read),                                                        //                                                .read
		.myCPU_data_master_readdata                                  (mycpu_data_master_readdata),                                                    //                                                .readdata
		.myCPU_data_master_readdatavalid                             (mycpu_data_master_readdatavalid),                                               //                                                .readdatavalid
		.myCPU_data_master_write                                     (mycpu_data_master_write),                                                       //                                                .write
		.myCPU_data_master_writedata                                 (mycpu_data_master_writedata),                                                   //                                                .writedata
		.myCPU_data_master_debugaccess                               (mycpu_data_master_debugaccess),                                                 //                                                .debugaccess
		.myCPU_instruction_master_address                            (mycpu_instruction_master_address),                                              //                        myCPU_instruction_master.address
		.myCPU_instruction_master_waitrequest                        (mycpu_instruction_master_waitrequest),                                          //                                                .waitrequest
		.myCPU_instruction_master_read                               (mycpu_instruction_master_read),                                                 //                                                .read
		.myCPU_instruction_master_readdata                           (mycpu_instruction_master_readdata),                                             //                                                .readdata
		.myCPU_instruction_master_readdatavalid                      (mycpu_instruction_master_readdatavalid),                                        //                                                .readdatavalid
		.audio_and_video_config_0_avalon_av_config_slave_address     (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address),     // audio_and_video_config_0_avalon_av_config_slave.address
		.audio_and_video_config_0_avalon_av_config_slave_write       (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write),       //                                                .write
		.audio_and_video_config_0_avalon_av_config_slave_read        (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read),        //                                                .read
		.audio_and_video_config_0_avalon_av_config_slave_readdata    (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata),    //                                                .readdata
		.audio_and_video_config_0_avalon_av_config_slave_writedata   (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata),   //                                                .writedata
		.audio_and_video_config_0_avalon_av_config_slave_byteenable  (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable),  //                                                .byteenable
		.audio_and_video_config_0_avalon_av_config_slave_waitrequest (mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest), //                                                .waitrequest
		.AudioCore_avalon_audio_slave_address                        (mm_interconnect_0_audiocore_avalon_audio_slave_address),                        //                    AudioCore_avalon_audio_slave.address
		.AudioCore_avalon_audio_slave_write                          (mm_interconnect_0_audiocore_avalon_audio_slave_write),                          //                                                .write
		.AudioCore_avalon_audio_slave_read                           (mm_interconnect_0_audiocore_avalon_audio_slave_read),                           //                                                .read
		.AudioCore_avalon_audio_slave_readdata                       (mm_interconnect_0_audiocore_avalon_audio_slave_readdata),                       //                                                .readdata
		.AudioCore_avalon_audio_slave_writedata                      (mm_interconnect_0_audiocore_avalon_audio_slave_writedata),                      //                                                .writedata
		.AudioCore_avalon_audio_slave_chipselect                     (mm_interconnect_0_audiocore_avalon_audio_slave_chipselect),                     //                                                .chipselect
		.GPIO_Expansion_s1_address                                   (mm_interconnect_0_gpio_expansion_s1_address),                                   //                               GPIO_Expansion_s1.address
		.GPIO_Expansion_s1_write                                     (mm_interconnect_0_gpio_expansion_s1_write),                                     //                                                .write
		.GPIO_Expansion_s1_readdata                                  (mm_interconnect_0_gpio_expansion_s1_readdata),                                  //                                                .readdata
		.GPIO_Expansion_s1_writedata                                 (mm_interconnect_0_gpio_expansion_s1_writedata),                                 //                                                .writedata
		.GPIO_Expansion_s1_chipselect                                (mm_interconnect_0_gpio_expansion_s1_chipselect),                                //                                                .chipselect
		.HEX0_s1_address                                             (mm_interconnect_0_hex0_s1_address),                                             //                                         HEX0_s1.address
		.HEX0_s1_write                                               (mm_interconnect_0_hex0_s1_write),                                               //                                                .write
		.HEX0_s1_readdata                                            (mm_interconnect_0_hex0_s1_readdata),                                            //                                                .readdata
		.HEX0_s1_writedata                                           (mm_interconnect_0_hex0_s1_writedata),                                           //                                                .writedata
		.HEX0_s1_chipselect                                          (mm_interconnect_0_hex0_s1_chipselect),                                          //                                                .chipselect
		.HEX1_s1_address                                             (mm_interconnect_0_hex1_s1_address),                                             //                                         HEX1_s1.address
		.HEX1_s1_write                                               (mm_interconnect_0_hex1_s1_write),                                               //                                                .write
		.HEX1_s1_readdata                                            (mm_interconnect_0_hex1_s1_readdata),                                            //                                                .readdata
		.HEX1_s1_writedata                                           (mm_interconnect_0_hex1_s1_writedata),                                           //                                                .writedata
		.HEX1_s1_chipselect                                          (mm_interconnect_0_hex1_s1_chipselect),                                          //                                                .chipselect
		.HEX2_s1_address                                             (mm_interconnect_0_hex2_s1_address),                                             //                                         HEX2_s1.address
		.HEX2_s1_write                                               (mm_interconnect_0_hex2_s1_write),                                               //                                                .write
		.HEX2_s1_readdata                                            (mm_interconnect_0_hex2_s1_readdata),                                            //                                                .readdata
		.HEX2_s1_writedata                                           (mm_interconnect_0_hex2_s1_writedata),                                           //                                                .writedata
		.HEX2_s1_chipselect                                          (mm_interconnect_0_hex2_s1_chipselect),                                          //                                                .chipselect
		.HEX3_s1_address                                             (mm_interconnect_0_hex3_s1_address),                                             //                                         HEX3_s1.address
		.HEX3_s1_write                                               (mm_interconnect_0_hex3_s1_write),                                               //                                                .write
		.HEX3_s1_readdata                                            (mm_interconnect_0_hex3_s1_readdata),                                            //                                                .readdata
		.HEX3_s1_writedata                                           (mm_interconnect_0_hex3_s1_writedata),                                           //                                                .writedata
		.HEX3_s1_chipselect                                          (mm_interconnect_0_hex3_s1_chipselect),                                          //                                                .chipselect
		.HEX4_s1_address                                             (mm_interconnect_0_hex4_s1_address),                                             //                                         HEX4_s1.address
		.HEX4_s1_write                                               (mm_interconnect_0_hex4_s1_write),                                               //                                                .write
		.HEX4_s1_readdata                                            (mm_interconnect_0_hex4_s1_readdata),                                            //                                                .readdata
		.HEX4_s1_writedata                                           (mm_interconnect_0_hex4_s1_writedata),                                           //                                                .writedata
		.HEX4_s1_chipselect                                          (mm_interconnect_0_hex4_s1_chipselect),                                          //                                                .chipselect
		.HEX5_s1_address                                             (mm_interconnect_0_hex5_s1_address),                                             //                                         HEX5_s1.address
		.HEX5_s1_write                                               (mm_interconnect_0_hex5_s1_write),                                               //                                                .write
		.HEX5_s1_readdata                                            (mm_interconnect_0_hex5_s1_readdata),                                            //                                                .readdata
		.HEX5_s1_writedata                                           (mm_interconnect_0_hex5_s1_writedata),                                           //                                                .writedata
		.HEX5_s1_chipselect                                          (mm_interconnect_0_hex5_s1_chipselect),                                          //                                                .chipselect
		.HEX6_s1_address                                             (mm_interconnect_0_hex6_s1_address),                                             //                                         HEX6_s1.address
		.HEX6_s1_write                                               (mm_interconnect_0_hex6_s1_write),                                               //                                                .write
		.HEX6_s1_readdata                                            (mm_interconnect_0_hex6_s1_readdata),                                            //                                                .readdata
		.HEX6_s1_writedata                                           (mm_interconnect_0_hex6_s1_writedata),                                           //                                                .writedata
		.HEX6_s1_chipselect                                          (mm_interconnect_0_hex6_s1_chipselect),                                          //                                                .chipselect
		.HEX7_s1_address                                             (mm_interconnect_0_hex7_s1_address),                                             //                                         HEX7_s1.address
		.HEX7_s1_write                                               (mm_interconnect_0_hex7_s1_write),                                               //                                                .write
		.HEX7_s1_readdata                                            (mm_interconnect_0_hex7_s1_readdata),                                            //                                                .readdata
		.HEX7_s1_writedata                                           (mm_interconnect_0_hex7_s1_writedata),                                           //                                                .writedata
		.HEX7_s1_chipselect                                          (mm_interconnect_0_hex7_s1_chipselect),                                          //                                                .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                       //                   jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                         //                                                .write
		.jtag_uart_0_avalon_jtag_slave_read                          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                          //                                                .read
		.jtag_uart_0_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                      //                                                .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                     //                                                .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                   //                                                .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                    //                                                .chipselect
		.KEYs_s1_address                                             (mm_interconnect_0_keys_s1_address),                                             //                                         KEYs_s1.address
		.KEYs_s1_write                                               (mm_interconnect_0_keys_s1_write),                                               //                                                .write
		.KEYs_s1_readdata                                            (mm_interconnect_0_keys_s1_readdata),                                            //                                                .readdata
		.KEYs_s1_writedata                                           (mm_interconnect_0_keys_s1_writedata),                                           //                                                .writedata
		.KEYs_s1_chipselect                                          (mm_interconnect_0_keys_s1_chipselect),                                          //                                                .chipselect
		.LEDG_s1_address                                             (mm_interconnect_0_ledg_s1_address),                                             //                                         LEDG_s1.address
		.LEDG_s1_write                                               (mm_interconnect_0_ledg_s1_write),                                               //                                                .write
		.LEDG_s1_readdata                                            (mm_interconnect_0_ledg_s1_readdata),                                            //                                                .readdata
		.LEDG_s1_writedata                                           (mm_interconnect_0_ledg_s1_writedata),                                           //                                                .writedata
		.LEDG_s1_chipselect                                          (mm_interconnect_0_ledg_s1_chipselect),                                          //                                                .chipselect
		.LEDR_s1_address                                             (mm_interconnect_0_ledr_s1_address),                                             //                                         LEDR_s1.address
		.LEDR_s1_write                                               (mm_interconnect_0_ledr_s1_write),                                               //                                                .write
		.LEDR_s1_readdata                                            (mm_interconnect_0_ledr_s1_readdata),                                            //                                                .readdata
		.LEDR_s1_writedata                                           (mm_interconnect_0_ledr_s1_writedata),                                           //                                                .writedata
		.LEDR_s1_chipselect                                          (mm_interconnect_0_ledr_s1_chipselect),                                          //                                                .chipselect
		.myCPU_jtag_debug_module_address                             (mm_interconnect_0_mycpu_jtag_debug_module_address),                             //                         myCPU_jtag_debug_module.address
		.myCPU_jtag_debug_module_write                               (mm_interconnect_0_mycpu_jtag_debug_module_write),                               //                                                .write
		.myCPU_jtag_debug_module_read                                (mm_interconnect_0_mycpu_jtag_debug_module_read),                                //                                                .read
		.myCPU_jtag_debug_module_readdata                            (mm_interconnect_0_mycpu_jtag_debug_module_readdata),                            //                                                .readdata
		.myCPU_jtag_debug_module_writedata                           (mm_interconnect_0_mycpu_jtag_debug_module_writedata),                           //                                                .writedata
		.myCPU_jtag_debug_module_byteenable                          (mm_interconnect_0_mycpu_jtag_debug_module_byteenable),                          //                                                .byteenable
		.myCPU_jtag_debug_module_waitrequest                         (mm_interconnect_0_mycpu_jtag_debug_module_waitrequest),                         //                                                .waitrequest
		.myCPU_jtag_debug_module_debugaccess                         (mm_interconnect_0_mycpu_jtag_debug_module_debugaccess),                         //                                                .debugaccess
		.sdram_s1_address                                            (mm_interconnect_0_sdram_s1_address),                                            //                                        sdram_s1.address
		.sdram_s1_write                                              (mm_interconnect_0_sdram_s1_write),                                              //                                                .write
		.sdram_s1_read                                               (mm_interconnect_0_sdram_s1_read),                                               //                                                .read
		.sdram_s1_readdata                                           (mm_interconnect_0_sdram_s1_readdata),                                           //                                                .readdata
		.sdram_s1_writedata                                          (mm_interconnect_0_sdram_s1_writedata),                                          //                                                .writedata
		.sdram_s1_byteenable                                         (mm_interconnect_0_sdram_s1_byteenable),                                         //                                                .byteenable
		.sdram_s1_readdatavalid                                      (mm_interconnect_0_sdram_s1_readdatavalid),                                      //                                                .readdatavalid
		.sdram_s1_waitrequest                                        (mm_interconnect_0_sdram_s1_waitrequest),                                        //                                                .waitrequest
		.sdram_s1_chipselect                                         (mm_interconnect_0_sdram_s1_chipselect),                                         //                                                .chipselect
		.switches_s1_address                                         (mm_interconnect_0_switches_s1_address),                                         //                                     switches_s1.address
		.switches_s1_write                                           (mm_interconnect_0_switches_s1_write),                                           //                                                .write
		.switches_s1_readdata                                        (mm_interconnect_0_switches_s1_readdata),                                        //                                                .readdata
		.switches_s1_writedata                                       (mm_interconnect_0_switches_s1_writedata),                                       //                                                .writedata
		.switches_s1_chipselect                                      (mm_interconnect_0_switches_s1_chipselect),                                      //                                                .chipselect
		.sysid_qsys_0_control_slave_address                          (mm_interconnect_0_sysid_qsys_0_control_slave_address),                          //                      sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                         (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                         //                                                .readdata
		.timer0_s1_address                                           (mm_interconnect_0_timer0_s1_address),                                           //                                       timer0_s1.address
		.timer0_s1_write                                             (mm_interconnect_0_timer0_s1_write),                                             //                                                .write
		.timer0_s1_readdata                                          (mm_interconnect_0_timer0_s1_readdata),                                          //                                                .readdata
		.timer0_s1_writedata                                         (mm_interconnect_0_timer0_s1_writedata),                                         //                                                .writedata
		.timer0_s1_chipselect                                        (mm_interconnect_0_timer0_s1_chipselect)                                         //                                                .chipselect
	);

	Nios2_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (mycpu_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (mycpu_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (clocks_reset_source_reset),           // reset_in1.reset
		.clk            (clocks_sys_clk_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
